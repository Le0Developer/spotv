module main

import sdl

// default dark theme of https://daisyui.com/theme-generator/
const background_100_color = sdl.Color{29, 35, 42, 255}
const background_200_color = sdl.Color{25, 30, 36, 255}
const background_300_color = sdl.Color{21, 25, 30, 255}
const text_color = sdl.Color{236, 249, 255, 255}
const muted_text_color = sdl.Color{136, 146, 161, 255}
const primary_color = sdl.Color{96, 93, 255, 255}
const primary_content_color = sdl.Color{237, 241, 254, 255}
const secondary_color = sdl.Color{244, 48, 152, 255}
const secondary_content_color = sdl.Color{249, 228, 240, 255}
const accent_color = sdl.Color{0, 211, 187, 255}
const accent_content_color = sdl.Color{8, 77, 73, 255}
const neutral_color = sdl.Color{9, 9, 11, 255}
const neutral_content_color = sdl.Color{228, 228, 231, 255}
const info_color = sdl.Color{0, 186, 254, 255}
const info_content_color = sdl.Color{4, 46, 73, 255}
const success_color = sdl.Color{0, 211, 144, 255}
const success_content_color = sdl.Color{0, 76, 57, 255}
const warning_color = sdl.Color{252, 183, 0, 255}
const warning_content_color = sdl.Color{121, 50, 5, 255}
const error_color = sdl.Color{255, 98, 125, 255}
const error_content_color = sdl.Color{77, 2, 24, 255}
