module main

#flag -framework Cocoa
#include <Cocoa/Cocoa.h>
#include "@DIR/window.m"

fn C.focusWindow()
fn C.setupWindow()
fn C.setupWindow2()
fn C.loseFocus()
